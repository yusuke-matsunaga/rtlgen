module ent1(
  input         port1,
  input         port2,
  input  [15:0] port3,
  output        oport
);
endmodule // ent1
